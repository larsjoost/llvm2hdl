library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity llvm_add is
  port (
    clk      : in  std_ulogic;
    sreset   : in  std_ulogic;
    s_tag    : in  std_ulogic_vector;
    s_tvalid : in  std_ulogic;
    s_tready : out std_ulogic;
    s_tdata  : in  std_ulogic_vector;
    m_tvalid : out std_ulogic;
    m_tready : in  std_ulogic;
    m_tag    : out std_ulogic_vector;
    m_tdata  : out std_ulogic_vector);
end entity llvm_add;

architecture rtl of llvm_add is

  constant data_width : positive := s_tdata'length/2;

  signal a_i, b_i, q_i : unsigned(0 to data_width - 1);

  signal s_tdata_i : std_ulogic_vector(0 to m_tdata'length - 1);
  
begin

  (a_i, b_i) <= unsigned(s_tdata);

  q_i <= a_i + b_i;

  s_tdata_i <= std_ulogic_vector(q_i);
  
  llvm_buffer_1 : entity work.llvm_buffer(rtl)
    port map (
      clk      => clk,
      sreset   => sreset,
      s_tag    => s_tag,
      s_tvalid => s_tvalid,
      s_tready => s_tready,
      s_tdata  => s_tdata_i,
      m_tvalid => m_tvalid,
      m_tready => m_tready,
      m_tag    => m_tag,
      m_tdata  => m_tdata);

end architecture rtl;
